// Created with Corsair v1.0.4

`ifndef __REGS_UFLASH_VH
`define __REGS_UFLASH_VH

`define UFLASH_BASE_ADDR 0
`define UFLASH_DATA_WIDTH 32
`define UFLASH_ADDR_WIDTH 32

// UFLASH_KEY1 - Unlock key for User Flash region
`define UFLASH_UFLASH_KEY1_ADDR 32'h0
`define UFLASH_UFLASH_KEY1_RESET 32'h0

// UFLASH_KEY1.KEY - 32-bit unlock key value(0x57494E44 - WIND)
`define UFLASH_UFLASH_KEY1_KEY_WIDTH 32
`define UFLASH_UFLASH_KEY1_KEY_LSB 0
`define UFLASH_UFLASH_KEY1_KEY_MASK 32'h0
`define UFLASH_UFLASH_KEY1_KEY_RESET 32'h0


// UFLASH_KEY2 - Unlock key for Text Flash region
`define UFLASH_UFLASH_KEY2_ADDR 32'h4
`define UFLASH_UFLASH_KEY2_RESET 32'h0

// UFLASH_KEY2.KEY - 32-bit unlock key value
`define UFLASH_UFLASH_KEY2_KEY_WIDTH 32
`define UFLASH_UFLASH_KEY2_KEY_LSB 0
`define UFLASH_UFLASH_KEY2_KEY_MASK 32'h4
`define UFLASH_UFLASH_KEY2_KEY_RESET 32'h0


// UFLASH_KEY3 - Unlock key for Boot Flash region
`define UFLASH_UFLASH_KEY3_ADDR 32'h8
`define UFLASH_UFLASH_KEY3_RESET 32'h0

// UFLASH_KEY3.KEY - 32-bit unlock key value
`define UFLASH_UFLASH_KEY3_KEY_WIDTH 32
`define UFLASH_UFLASH_KEY3_KEY_LSB 0
`define UFLASH_UFLASH_KEY3_KEY_MASK 32'h8
`define UFLASH_UFLASH_KEY3_KEY_RESET 32'h0


// UFLASH_CR - Flash Control Register
`define UFLASH_UFLASH_CR_ADDR 32'hc
`define UFLASH_UFLASH_CR_RESET 32'h0

// UFLASH_CR.USER_EN - Enable access to User region
`define UFLASH_UFLASH_CR_USER_EN_WIDTH 1
`define UFLASH_UFLASH_CR_USER_EN_LSB 0
`define UFLASH_UFLASH_CR_USER_EN_MASK 32'hc
`define UFLASH_UFLASH_CR_USER_EN_RESET 1'h0

// UFLASH_CR.TEXT_EN - Enable access to Text region
`define UFLASH_UFLASH_CR_TEXT_EN_WIDTH 1
`define UFLASH_UFLASH_CR_TEXT_EN_LSB 1
`define UFLASH_UFLASH_CR_TEXT_EN_MASK 32'hc
`define UFLASH_UFLASH_CR_TEXT_EN_RESET 1'h0

// UFLASH_CR.BOOT_EN - Enable access to Boot region
`define UFLASH_UFLASH_CR_BOOT_EN_WIDTH 1
`define UFLASH_UFLASH_CR_BOOT_EN_LSB 2
`define UFLASH_UFLASH_CR_BOOT_EN_MASK 32'hc
`define UFLASH_UFLASH_CR_BOOT_EN_RESET 1'h0

// UFLASH_CR.PROG_EN - Program enable
`define UFLASH_UFLASH_CR_PROG_EN_WIDTH 1
`define UFLASH_UFLASH_CR_PROG_EN_LSB 3
`define UFLASH_UFLASH_CR_PROG_EN_MASK 32'hc
`define UFLASH_UFLASH_CR_PROG_EN_RESET 1'h0

// UFLASH_CR.READ_EN - Read enable
`define UFLASH_UFLASH_CR_READ_EN_WIDTH 1
`define UFLASH_UFLASH_CR_READ_EN_LSB 4
`define UFLASH_UFLASH_CR_READ_EN_MASK 32'hc
`define UFLASH_UFLASH_CR_READ_EN_RESET 1'h0

// UFLASH_CR.ERASE_EN - Erase enable
`define UFLASH_UFLASH_CR_ERASE_EN_WIDTH 1
`define UFLASH_UFLASH_CR_ERASE_EN_LSB 5
`define UFLASH_UFLASH_CR_ERASE_EN_MASK 32'hc
`define UFLASH_UFLASH_CR_ERASE_EN_RESET 1'h0

// UFLASH_CR.MODE - Flash operation mode
`define UFLASH_UFLASH_CR_MODE_WIDTH 2
`define UFLASH_UFLASH_CR_MODE_LSB 6
`define UFLASH_UFLASH_CR_MODE_MASK 32'hc
`define UFLASH_UFLASH_CR_MODE_RESET 2'h0
`define UFLASH_UFLASH_CR_MODE_READ 2'h0 //Read mode
`define UFLASH_UFLASH_CR_MODE_PROGRAM 2'h1 //Program mode
`define UFLASH_UFLASH_CR_MODE_ERASE 2'h2 //Erase mode
`define UFLASH_UFLASH_CR_MODE_IDLE 2'h3 //Idle mode


// UFLASH_SR - Flash Status Register
`define UFLASH_UFLASH_SR_ADDR 32'h10
`define UFLASH_UFLASH_SR_RESET 32'h0

// UFLASH_SR.ERRA_USER - Error unauthorized access to User region
`define UFLASH_UFLASH_SR_ERRA_USER_WIDTH 1
`define UFLASH_UFLASH_SR_ERRA_USER_LSB 0
`define UFLASH_UFLASH_SR_ERRA_USER_MASK 32'h10
`define UFLASH_UFLASH_SR_ERRA_USER_RESET 1'h0

// UFLASH_SR.ERRA_TEXT - Error unauthorized access to Text region
`define UFLASH_UFLASH_SR_ERRA_TEXT_WIDTH 1
`define UFLASH_UFLASH_SR_ERRA_TEXT_LSB 1
`define UFLASH_UFLASH_SR_ERRA_TEXT_MASK 32'h10
`define UFLASH_UFLASH_SR_ERRA_TEXT_RESET 1'h0

// UFLASH_SR.ERRA_BOOT - Error unauthorized access to Boot region
`define UFLASH_UFLASH_SR_ERRA_BOOT_WIDTH 1
`define UFLASH_UFLASH_SR_ERRA_BOOT_LSB 2
`define UFLASH_UFLASH_SR_ERRA_BOOT_MASK 32'h10
`define UFLASH_UFLASH_SR_ERRA_BOOT_RESET 1'h0

// UFLASH_SR.ERRA_OVF - Error address overflow
`define UFLASH_UFLASH_SR_ERRA_OVF_WIDTH 1
`define UFLASH_UFLASH_SR_ERRA_OVF_LSB 3
`define UFLASH_UFLASH_SR_ERRA_OVF_MASK 32'h10
`define UFLASH_UFLASH_SR_ERRA_OVF_RESET 1'h0

// UFLASH_SR.RD_DONE - Read operation finished
`define UFLASH_UFLASH_SR_RD_DONE_WIDTH 1
`define UFLASH_UFLASH_SR_RD_DONE_LSB 4
`define UFLASH_UFLASH_SR_RD_DONE_MASK 32'h10
`define UFLASH_UFLASH_SR_RD_DONE_RESET 1'h0

// UFLASH_SR.PROG_DONE - Program operation finished
`define UFLASH_UFLASH_SR_PROG_DONE_WIDTH 1
`define UFLASH_UFLASH_SR_PROG_DONE_LSB 5
`define UFLASH_UFLASH_SR_PROG_DONE_MASK 32'h10
`define UFLASH_UFLASH_SR_PROG_DONE_RESET 1'h0

// UFLASH_SR.ERASE_DONE - Erase operation finished
`define UFLASH_UFLASH_SR_ERASE_DONE_WIDTH 1
`define UFLASH_UFLASH_SR_ERASE_DONE_LSB 6
`define UFLASH_UFLASH_SR_ERASE_DONE_MASK 32'h10
`define UFLASH_UFLASH_SR_ERASE_DONE_RESET 1'h0


// UFLASH_XADR - Flash X Address Register
`define UFLASH_UFLASH_XADR_ADDR 32'h14
`define UFLASH_UFLASH_XADR_RESET 32'h0

// UFLASH_XADR.XADR - Flash X address (row / page select)
`define UFLASH_UFLASH_XADR_XADR_WIDTH 16
`define UFLASH_UFLASH_XADR_XADR_LSB 0
`define UFLASH_UFLASH_XADR_XADR_MASK 32'h14
`define UFLASH_UFLASH_XADR_XADR_RESET 16'h0


// UFLASH_YADR - Flash Y Address Register
`define UFLASH_UFLASH_YADR_ADDR 32'h18
`define UFLASH_UFLASH_YADR_RESET 32'h0

// UFLASH_YADR.YADR - Flash Y address (column / word select)
`define UFLASH_UFLASH_YADR_YADR_WIDTH 8
`define UFLASH_UFLASH_YADR_YADR_LSB 0
`define UFLASH_UFLASH_YADR_YADR_MASK 32'h18
`define UFLASH_UFLASH_YADR_YADR_RESET 8'h0


// UFLASH_DOR - Flash data out Register
`define UFLASH_UFLASH_DOR_ADDR 32'h1c
`define UFLASH_UFLASH_DOR_RESET 32'h0

// UFLASH_DOR.DO - 32BIT READ DATA
`define UFLASH_UFLASH_DOR_DO_WIDTH 32
`define UFLASH_UFLASH_DOR_DO_LSB 0
`define UFLASH_UFLASH_DOR_DO_MASK 32'h1c
`define UFLASH_UFLASH_DOR_DO_RESET 32'h0


// UFLASH_DIR - Flash data in Register
`define UFLASH_UFLASH_DIR_ADDR 32'h20
`define UFLASH_UFLASH_DIR_RESET 32'h0

// UFLASH_DIR.DI - 32BIT PROGRAM DATA
`define UFLASH_UFLASH_DIR_DI_WIDTH 32
`define UFLASH_UFLASH_DIR_DI_LSB 0
`define UFLASH_UFLASH_DIR_DI_MASK 32'h20
`define UFLASH_UFLASH_DIR_DI_RESET 32'h0


`endif // __REGS_UFLASH_VH