// Created with Corsair v1.0.4

`ifndef __REGS_GPIO_VH
`define __REGS_GPIO_VH

`define GPIO_BASE_ADDR 1073741824
`define GPIO_DATA_WIDTH 32
`define GPIO_ADDR_WIDTH 32

// GPIO_IO - GPIO Read/Write Register
`define GPIO_GPIO_IO_ADDR 32'h0
`define GPIO_GPIO_IO_RESET 32'h0

// GPIO_IO.GPIO_0 - GPIO0
`define GPIO_GPIO_IO_GPIO_0_WIDTH 1
`define GPIO_GPIO_IO_GPIO_0_LSB 0
`define GPIO_GPIO_IO_GPIO_0_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_0_RESET 1'h0

// GPIO_IO.GPIO_1 - GPIO1
`define GPIO_GPIO_IO_GPIO_1_WIDTH 1
`define GPIO_GPIO_IO_GPIO_1_LSB 1
`define GPIO_GPIO_IO_GPIO_1_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_1_RESET 1'h0

// GPIO_IO.GPIO_2 - GPIO2
`define GPIO_GPIO_IO_GPIO_2_WIDTH 1
`define GPIO_GPIO_IO_GPIO_2_LSB 2
`define GPIO_GPIO_IO_GPIO_2_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_2_RESET 1'h0

// GPIO_IO.GPIO_3 - GPIO3
`define GPIO_GPIO_IO_GPIO_3_WIDTH 1
`define GPIO_GPIO_IO_GPIO_3_LSB 3
`define GPIO_GPIO_IO_GPIO_3_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_3_RESET 1'h0

// GPIO_IO.GPIO_4 - GPIO4
`define GPIO_GPIO_IO_GPIO_4_WIDTH 1
`define GPIO_GPIO_IO_GPIO_4_LSB 4
`define GPIO_GPIO_IO_GPIO_4_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_4_RESET 1'h0

// GPIO_IO.GPIO_5 - GPIO5
`define GPIO_GPIO_IO_GPIO_5_WIDTH 1
`define GPIO_GPIO_IO_GPIO_5_LSB 5
`define GPIO_GPIO_IO_GPIO_5_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_5_RESET 1'h0

// GPIO_IO.GPIO_6 - GPIO6
`define GPIO_GPIO_IO_GPIO_6_WIDTH 1
`define GPIO_GPIO_IO_GPIO_6_LSB 6
`define GPIO_GPIO_IO_GPIO_6_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_6_RESET 1'h0

// GPIO_IO.GPIO_7 - GPIO7
`define GPIO_GPIO_IO_GPIO_7_WIDTH 1
`define GPIO_GPIO_IO_GPIO_7_LSB 7
`define GPIO_GPIO_IO_GPIO_7_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_7_RESET 1'h0

// GPIO_IO.GPIO_8 - GPIO8
`define GPIO_GPIO_IO_GPIO_8_WIDTH 1
`define GPIO_GPIO_IO_GPIO_8_LSB 8
`define GPIO_GPIO_IO_GPIO_8_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_8_RESET 1'h0

// GPIO_IO.GPIO_9 - GPIO9
`define GPIO_GPIO_IO_GPIO_9_WIDTH 1
`define GPIO_GPIO_IO_GPIO_9_LSB 9
`define GPIO_GPIO_IO_GPIO_9_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_9_RESET 1'h0

// GPIO_IO.GPIO_10 - GPIO10
`define GPIO_GPIO_IO_GPIO_10_WIDTH 1
`define GPIO_GPIO_IO_GPIO_10_LSB 10
`define GPIO_GPIO_IO_GPIO_10_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_10_RESET 1'h0

// GPIO_IO.GPIO_11 - GPIO11
`define GPIO_GPIO_IO_GPIO_11_WIDTH 1
`define GPIO_GPIO_IO_GPIO_11_LSB 11
`define GPIO_GPIO_IO_GPIO_11_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_11_RESET 1'h0

// GPIO_IO.GPIO_12 - GPIO12
`define GPIO_GPIO_IO_GPIO_12_WIDTH 1
`define GPIO_GPIO_IO_GPIO_12_LSB 12
`define GPIO_GPIO_IO_GPIO_12_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_12_RESET 1'h0

// GPIO_IO.GPIO_13 - GPIO13
`define GPIO_GPIO_IO_GPIO_13_WIDTH 1
`define GPIO_GPIO_IO_GPIO_13_LSB 13
`define GPIO_GPIO_IO_GPIO_13_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_13_RESET 1'h0

// GPIO_IO.GPIO_14 - GPIO14
`define GPIO_GPIO_IO_GPIO_14_WIDTH 1
`define GPIO_GPIO_IO_GPIO_14_LSB 14
`define GPIO_GPIO_IO_GPIO_14_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_14_RESET 1'h0

// GPIO_IO.GPIO_15 - GPIO15
`define GPIO_GPIO_IO_GPIO_15_WIDTH 1
`define GPIO_GPIO_IO_GPIO_15_LSB 15
`define GPIO_GPIO_IO_GPIO_15_MASK 32'h0
`define GPIO_GPIO_IO_GPIO_15_RESET 1'h0


// GPIO_config - GPIO config Register 0 output, 1 input
`define GPIO_GPIO_CONFIG_ADDR 32'h4
`define GPIO_GPIO_CONFIG_RESET 32'h0

// GPIO_config.GPIO_0config - GPIO0_config
`define GPIO_GPIO_CONFIG_GPIO_0CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_0CONFIG_LSB 0
`define GPIO_GPIO_CONFIG_GPIO_0CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_0CONFIG_RESET 1'h0

// GPIO_config.GPIO_1config - GPIO1_config
`define GPIO_GPIO_CONFIG_GPIO_1CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_1CONFIG_LSB 1
`define GPIO_GPIO_CONFIG_GPIO_1CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_1CONFIG_RESET 1'h0

// GPIO_config.GPIO_2config - GPIO2_config
`define GPIO_GPIO_CONFIG_GPIO_2CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_2CONFIG_LSB 2
`define GPIO_GPIO_CONFIG_GPIO_2CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_2CONFIG_RESET 1'h0

// GPIO_config.GPIO_3config - GPIO3_config
`define GPIO_GPIO_CONFIG_GPIO_3CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_3CONFIG_LSB 3
`define GPIO_GPIO_CONFIG_GPIO_3CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_3CONFIG_RESET 1'h0

// GPIO_config.GPIO_4config - GPIO4_config
`define GPIO_GPIO_CONFIG_GPIO_4CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_4CONFIG_LSB 4
`define GPIO_GPIO_CONFIG_GPIO_4CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_4CONFIG_RESET 1'h0

// GPIO_config.GPIO_5config - GPIO5_config
`define GPIO_GPIO_CONFIG_GPIO_5CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_5CONFIG_LSB 5
`define GPIO_GPIO_CONFIG_GPIO_5CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_5CONFIG_RESET 1'h0

// GPIO_config.GPIO_6config - GPIO6_config
`define GPIO_GPIO_CONFIG_GPIO_6CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_6CONFIG_LSB 6
`define GPIO_GPIO_CONFIG_GPIO_6CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_6CONFIG_RESET 1'h0

// GPIO_config.GPIO_7config - GPIO7_config
`define GPIO_GPIO_CONFIG_GPIO_7CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_7CONFIG_LSB 7
`define GPIO_GPIO_CONFIG_GPIO_7CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_7CONFIG_RESET 1'h0

// GPIO_config.GPIO_8config - GPIO8_config
`define GPIO_GPIO_CONFIG_GPIO_8CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_8CONFIG_LSB 8
`define GPIO_GPIO_CONFIG_GPIO_8CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_8CONFIG_RESET 1'h0

// GPIO_config.GPIO_9config - GPIO9_config
`define GPIO_GPIO_CONFIG_GPIO_9CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_9CONFIG_LSB 9
`define GPIO_GPIO_CONFIG_GPIO_9CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_9CONFIG_RESET 1'h0

// GPIO_config.GPIO_10config - GPIO10_config
`define GPIO_GPIO_CONFIG_GPIO_10CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_10CONFIG_LSB 10
`define GPIO_GPIO_CONFIG_GPIO_10CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_10CONFIG_RESET 1'h0

// GPIO_config.GPIO_11config - GPIO11_config
`define GPIO_GPIO_CONFIG_GPIO_11CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_11CONFIG_LSB 11
`define GPIO_GPIO_CONFIG_GPIO_11CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_11CONFIG_RESET 1'h0

// GPIO_config.GPIO_12config - GPIO12_config
`define GPIO_GPIO_CONFIG_GPIO_12CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_12CONFIG_LSB 12
`define GPIO_GPIO_CONFIG_GPIO_12CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_12CONFIG_RESET 1'h0

// GPIO_config.GPIO_13config - GPIO13_config
`define GPIO_GPIO_CONFIG_GPIO_13CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_13CONFIG_LSB 13
`define GPIO_GPIO_CONFIG_GPIO_13CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_13CONFIG_RESET 1'h0

// GPIO_config.GPIO_14config - GPIO14_config
`define GPIO_GPIO_CONFIG_GPIO_14CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_14CONFIG_LSB 14
`define GPIO_GPIO_CONFIG_GPIO_14CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_14CONFIG_RESET 1'h0

// GPIO_config.GPIO_15config - GPIO15_config
`define GPIO_GPIO_CONFIG_GPIO_15CONFIG_WIDTH 1
`define GPIO_GPIO_CONFIG_GPIO_15CONFIG_LSB 15
`define GPIO_GPIO_CONFIG_GPIO_15CONFIG_MASK 32'h4
`define GPIO_GPIO_CONFIG_GPIO_15CONFIG_RESET 1'h0


`endif // __REGS_GPIO_VH