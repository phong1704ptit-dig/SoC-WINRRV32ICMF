//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Wed Sep 17 13:03:05 2025

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [31:0] douta;
output [31:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [11:0] ada;
input [31:0] dina;
input [11:0] adb;
input [31:0] dinb;

wire [11:0] dpb_inst_0_douta_w;
wire [11:0] dpb_inst_0_doutb_w;
wire [11:0] dpb_inst_1_douta_w;
wire [11:0] dpb_inst_1_doutb_w;
wire [11:0] dpb_inst_2_douta_w;
wire [11:0] dpb_inst_2_doutb_w;
wire [11:0] dpb_inst_3_douta_w;
wire [11:0] dpb_inst_3_doutb_w;
wire [11:0] dpb_inst_4_douta_w;
wire [11:0] dpb_inst_4_doutb_w;
wire [11:0] dpb_inst_5_douta_w;
wire [11:0] dpb_inst_5_doutb_w;
wire [11:0] dpb_inst_6_douta_w;
wire [11:0] dpb_inst_6_doutb_w;
wire [11:0] dpb_inst_7_douta_w;
wire [11:0] dpb_inst_7_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[11:0],douta[3:0]}),
    .DOB({dpb_inst_0_doutb_w[11:0],doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 4;
defparam dpb_inst_0.BIT_WIDTH_1 = 4;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h37733333333FF33333373337333733337733333333333333333F3F3333333F37;
defparam dpb_inst_0.INIT_RAM_01 = 256'h3337333737373373373333F33373733373773337373337373333337333733373;
defparam dpb_inst_0.INIT_RAM_02 = 256'h733333333337333333333333333333333333333333333333333333F337733F33;
defparam dpb_inst_0.INIT_RAM_03 = 256'h333F3337F3F33F33F33F33F33F333F333F333F333F333F333733333333FFFFF3;
defparam dpb_inst_0.INIT_RAM_04 = 256'h33333333333333FF3F333333333333333333333337333333333733333333333F;
defparam dpb_inst_0.INIT_RAM_05 = 256'h3333333333333337773333733733373333733333333333337733333F3F33F333;
defparam dpb_inst_0.INIT_RAM_06 = 256'h733F33F333333333333333333333333F33333333333333333373373773373333;
defparam dpb_inst_0.INIT_RAM_07 = 256'h3733F3333733F333373333333333FF37333FF337733333333F37F333F37F33F3;
defparam dpb_inst_0.INIT_RAM_08 = 256'h3733373337333733373FFFF3333FF373373733333333F37F333F37F33F3733F3;
defparam dpb_inst_0.INIT_RAM_09 = 256'hF333F3333F333333333333333333333373333733333333333333FF3F33F33733;
defparam dpb_inst_0.INIT_RAM_0A = 256'h33333733F3F33F333773333333333333333333333333F333F333F33333333333;
defparam dpb_inst_0.INIT_RAM_0B = 256'h333333F3337F33333333333F333F333F33333333333F333F3333F33333333333;
defparam dpb_inst_0.INIT_RAM_0C = 256'h33373F3F33F33F33F333333333333F333F333F33333333333F333F333F333333;
defparam dpb_inst_0.INIT_RAM_0D = 256'h3F333F333F33333333333F333F333F33333333333333F3337F33333333333373;
defparam dpb_inst_0.INIT_RAM_0E = 256'h3333333F33F33F33F33333333333373333F333F333F3333F3333333333333333;
defparam dpb_inst_0.INIT_RAM_0F = 256'h333F3F333333333333333F333F33F33333333333333333333733373333333333;
defparam dpb_inst_0.INIT_RAM_10 = 256'h3F3333333333333333333333733F33377333333333333333333333333333333F;
defparam dpb_inst_0.INIT_RAM_11 = 256'h3333333333F333F33F333333333333333333F333F3F333333333333333F333F3;
defparam dpb_inst_0.INIT_RAM_12 = 256'h3333333333333F3337F33333333333333337333373F3337F3333F333F3F33333;
defparam dpb_inst_0.INIT_RAM_13 = 256'h3F333F3333F3333F33333333333333333F333F333F33333333333F333F333F33;
defparam dpb_inst_0.INIT_RAM_14 = 256'h373333333333333333333733333333F33F33F333333333333333333333337333;
defparam dpb_inst_0.INIT_RAM_15 = 256'h000000000000000000000000000000000000000073F33373F33373F33F33373F;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[11:0],douta[7:4]}),
    .DOB({dpb_inst_1_doutb_w[11:0],doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b1;
defparam dpb_inst_1.READ_MODE1 = 1'b1;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 4;
defparam dpb_inst_1.BIT_WIDTH_1 = 4;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h8B61088E0B9E691222162983E98B2102B610811E80298E902986262212217E11;
defparam dpb_inst_1.INIT_RAM_01 = 256'hBB9B81130B2B68B2161882E2B138B22162B62B9B2B169B0B692B313099B29839;
defparam dpb_inst_1.INIT_RAM_02 = 256'h39961619998BE1971808080808080880886F222222222222222221621B618E12;
defparam dpb_inst_1.INIT_RAM_03 = 256'h129E129369E12E12E12E12E12E129E121E129E121E129E121B222222216E6E62;
defparam dpb_inst_1.INIT_RAM_04 = 256'h96BEE8B191B13B6E1699282222222220808008009B912226B21610808088E99E;
defparam dpb_inst_1.INIT_RAM_05 = 256'h2102021020202983B67979B796239B0239B0210210210210B61880869E116169;
defparam dpb_inst_1.INIT_RAM_06 = 256'h391E91EB19199B3B393193B3B1B9991E919191912222226B2162BB83620B2020;
defparam dpb_inst_1.INIT_RAM_07 = 256'h1391E9191391E9191319222222216E13E966E113618080808E13E916E13E91E1;
defparam dpb_inst_1.INIT_RAM_08 = 256'h23F22B722BF22B722BFEEEE22216E13E9B6610808088E13E916E13E91E1391E9;
defparam dpb_inst_1.INIT_RAM_09 = 256'hE191E1199E1991B3BB3361B8BB11161136999B692222222222216E1E08E22BF2;
defparam dpb_inst_1.INIT_RAM_0A = 256'hB1116361696B161E1B610198080880808B9966B6B919E199E199E193166B6B91;
defparam dpb_inst_1.INIT_RAM_0B = 256'hBB13B361E1B6B9966B6B919E191E199E193166B6B91E199E1191E11991361B8B;
defparam dpb_inst_1.INIT_RAM_0C = 256'h116B6696B16B96B16331966B6B919E199E199E193166B6B91E199E119E9B1993;
defparam dpb_inst_1.INIT_RAM_0D = 256'h9E191E119E19B16636311E191E119E1B1913BB9BBBB361E1B61BB9B6B18B93B1;
defparam dpb_inst_1.INIT_RAM_0E = 256'h22222216916B163169EEB3191631336B39E191E191E9111E9B1B1111166B6B91;
defparam dpb_inst_1.INIT_RAM_0F = 256'h199E9E193B33393BB6B91E191E99E19913BBBB631B8BB11163699B6912222222;
defparam dpb_inst_1.INIT_RAM_10 = 256'h1E119339BBBB633B98BB111636161E1B6180808080808089333BBB1B3363119E;
defparam dpb_inst_1.INIT_RAM_11 = 256'h3393BB6B91E191E99E1991BB33393BB6B919E191E9E19B3BBB9BB36311E199E9;
defparam dpb_inst_1.INIT_RAM_12 = 256'h311B93B93BBBB61E1B691BBB1B666390B93B1116BE61E1B63111E199E9E193B3;
defparam dpb_inst_1.INIT_RAM_13 = 256'hBE191E1999E9111E91191331166B6B919E119E119E19B166B6B91E191E119E1B;
defparam dpb_inst_1.INIT_RAM_14 = 256'h96E193B61E916696191666E19369116B16B16B3B3BBBB39BBB666B319193B6B9;
defparam dpb_inst_1.INIT_RAM_15 = 256'h000000000000000000000000000000000000000063E3EB61E66963E9B6B6361E;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[11:0],douta[11:8]}),
    .DOB({dpb_inst_2_doutb_w[11:0],doutb[11:8]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[11:8]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[11:8]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b1;
defparam dpb_inst_2.READ_MODE1 = 1'b1;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 4;
defparam dpb_inst_2.BIT_WIDTH_1 = 4;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'h670194085740049246100777A777077470140006776776774770406E44610011;
defparam dpb_inst_2.INIT_RAM_01 = 256'h7766777677076776101404007557446104700777476277772707766777527776;
defparam dpb_inst_2.INIT_RAM_02 = 256'h77707077747767701FFEE88776655433208768ACE02468ACE024610077010050;
defparam dpb_inst_2.INIT_RAM_03 = 256'h50705079040500500500500500507050B050A050A0509050942468ACE1000002;
defparam dpb_inst_2.INIT_RAM_04 = 256'h9C7CE77775497700506967420ECA86476655883E77498ACE7E101BAA9940A740;
defparam dpb_inst_2.INIT_RAM_05 = 256'h2772727727260667700707707007667076670770770770777010994060550507;
defparam dpb_inst_2.INIT_RAM_06 = 256'h54906605566757775777676777667AB05566994A2468ACE7E102767700774747;
defparam dpb_inst_2.INIT_RAM_07 = 256'h664B0556669A055666942468ACE1005547600555010BAA994055055A05505505;
defparam dpb_inst_2.INIT_RAM_08 = 256'hC9720766476A875EC75000024610055C77801BAA99400550550055055055A906;
defparam dpb_inst_2.INIT_RAM_09 = 256'h05540595B05B5B4C97C7E777767778CA7474974A2468CE0246A10050550A847E;
defparam dpb_inst_2.INIT_RAM_0A = 256'h677747C70A06907C7601A55CCBBA9944077A644A4454055B05A505549A46A665;
defparam dpb_inst_2.INIT_RAM_0B = 256'h75B49707076077B244A4454055B05B505549646A665055B0595B05B5AA4C7777;
defparam dpb_inst_2.INIT_RAM_0C = 256'h774760B06907A0690A49A247A7757055B05A505549646A665055A05950B455BA;
defparam dpb_inst_2.INIT_RAM_0D = 256'h7055C059505544E47A775055905450C955CA57C4B6BB070770A767787B777577;
defparam dpb_inst_2.INIT_RAM_0E = 256'h468EAC107A07907407026786806657667605530557055580575853439A47A775;
defparam dpb_inst_2.INIT_RAM_0F = 256'h55A05055B777767672775055B05A05A5A44975C977776777270797A4468ACE02;
defparam dpb_inst_2.INIT_RAM_10 = 256'hB05B54AA57B9E974767677727C70727601DDCCBBAA9944055557777775255570;
defparam dpb_inst_2.INIT_RAM_11 = 256'h7767672775055B05A05A5A47777676727757055B050554777767672775055405;
defparam dpb_inst_2.INIT_RAM_12 = 256'h95D4597CBBB6A0787705544644C40AAA7787777C760727605454055A05055B77;
defparam dpb_inst_2.INIT_RAM_13 = 256'h705530557505558055455474B245A555505C505B5055D4647A775055C05450D9;
defparam dpb_inst_2.INIT_RAM_14 = 256'h206665565A668A6C5566006655465605B0740557A545757669CE675878656676;
defparam dpb_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000050585050CA2050250585050;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[11:0],douta[15:12]}),
    .DOB({dpb_inst_3_doutb_w[11:0],doutb[15:12]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[15:12]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[15:12]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b1;
defparam dpb_inst_3.READ_MODE1 = 1'b1;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 4;
defparam dpb_inst_3.BIT_WIDTH_1 = 4;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'hA0802221C08F000222082F209FA0A6AA0802200422282D022820202202200004;
defparam dpb_inst_3.INIT_RAM_01 = 256'hEF8C2170A1A18A1208022AF8000A12208A188880A10C81A180A670CA9F02821F;
defparam dpb_inst_3.INIT_RAM_02 = 256'h0D98080D98A090F0022222222222222222C2222222222222222220FA01802F02;
defparam dpb_inst_3.INIT_RAM_03 = 256'h020F020000F0AF0AF0AF0AF0AF0A0F0A0F0A0F0A0F0A0F0A0022222220FFFFF2;
defparam dpb_inst_3.INIT_RAM_04 = 256'h89E79A809088300F00002A222222222AAAAAAAAA80802228620802222222D08F;
defparam dpb_inst_3.INIT_RAM_05 = 256'hA6AAAA6AAA2220220890981908A682AA780AA6AA7AA6AA7A0802222F0F70F0C0;
defparam dpb_inst_3.INIT_RAM_06 = 256'h08000008108958038981D08B0981D800080880802222228E2082E8208AA0AAAA;
defparam dpb_inst_3.INIT_RAM_07 = 256'h0280080004800880048022222220FF00E09FF000802222222F00F808F00F80F0;
defparam dpb_inst_3.INIT_RAM_08 = 256'h212AA12AA12AA12AA12FFFF2220FF00E889802222222F00F808F00F80F008000;
defparam dpb_inst_3.INIT_RAM_09 = 256'h00000800D0090D9E1D90808C851337880F800090222222222220FF0FA2FAA122;
defparam dpb_inst_3.INIT_RAM_0A = 256'h51337000F8F80F0700802802222222222E18FF8FED190000080000080FF8FED1;
defparam dpb_inst_3.INIT_RAM_0B = 256'hD9DD10F0700FE18FF8FED190080000000880FF8FED10080000050098D08908C8;
defparam dpb_inst_3.INIT_RAM_0C = 256'h3BF0EF8F80F88F80F6818FF8FED110000080000080FF8FE51000008000D9009E;
defparam dpb_inst_3.INIT_RAM_0D = 256'h10880000008800778765108800000051889E9DDDE950F0F00F0EBBB980C88D01;
defparam dpb_inst_3.INIT_RAM_0E = 256'h2222220F00F80F00F89789591E0D00F8050DD00D000D5100065815190FF8FED1;
defparam dpb_inst_3.INIT_RAM_0F = 256'h0000800080707BBB8FE51080008D0890D1E1598008C8513370F8009802222222;
defparam dpb_inst_3.INIT_RAM_10 = 256'h508981ED95D108880C851337000F07008022222222222220508F0F3338765110;
defparam dpb_inst_3.INIT_RAM_11 = 256'h07BBB8FE51080008D0890D80707BBB8FED1108800008808F0FB3387651088000;
defparam dpb_inst_3.INIT_RAM_12 = 256'h6091859DDE598F0F00F8083880F7100C88D013BF0EF0700F6511000008000807;
defparam dpb_inst_3.INIT_RAM_13 = 256'h800D000D090D5100D55916810FF8FED110808000008880FF8FE5100800000051;
defparam dpb_inst_3.INIT_RAM_14 = 256'h8895D68E06915700008C4891D08F00F80F80FD6D98B08088B81F688591D00F85;
defparam dpb_inst_3.INIT_RAM_15 = 256'h000000000000000000000000000000000000000080F05088F4C880F80F04088F;

DPB dpb_inst_4 (
    .DOA({dpb_inst_4_douta_w[11:0],douta[19:16]}),
    .DOB({dpb_inst_4_doutb_w[11:0],doutb[19:16]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[19:16]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[19:16]})
);

defparam dpb_inst_4.READ_MODE0 = 1'b1;
defparam dpb_inst_4.READ_MODE1 = 1'b1;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 4;
defparam dpb_inst_4.BIT_WIDTH_1 = 4;
defparam dpb_inst_4.BLK_SEL_0 = 3'b000;
defparam dpb_inst_4.BLK_SEL_1 = 3'b000;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'h70011115794F0051111077707770777700111007444747044740404411110010;
defparam dpb_inst_4.INIT_RAM_01 = 256'h776F677070707701101114F7550401110700777070777070605776F577077706;
defparam dpb_inst_4.INIT_RAM_02 = 256'h074707077770707011111111111111111170111111111111111111F700011F06;
defparam dpb_inst_4.INIT_RAM_03 = 256'h090F090000F04F04F04F04F04F040F040F040F040F040F040011111111FFFFF7;
defparam dpb_inst_4.INIT_RAM_04 = 256'h976947719547990F00001711111111177777777770551117511011111111704F;
defparam dpb_inst_4.INIT_RAM_05 = 256'h7777777777777070007077070077607776F77777777777770011111F0F55F070;
defparam dpb_inst_4.INIT_RAM_06 = 256'h055000055997577577677767747A4550A5966655111111761107707007707777;
defparam dpb_inst_4.INIT_RAM_07 = 256'h605504906F5504506F5511111111FF50704FF550011111111F50F494F50FABF5;
defparam dpb_inst_4.INIT_RAM_08 = 256'h9007700770077007700FFFF1111FF507714011111111F50FA94F50F9AF505500;
defparam dpb_inst_4.INIT_RAM_09 = 256'h0CB50B55B0C9B9A76A5770777677665615756065111111111111FF0F49F44009;
defparam dpb_inst_4.INIT_RAM_0A = 256'h67766160FAF69F06000117A111111111179A4494445404B50B5504B696696645;
defparam dpb_inst_4.INIT_RAM_0B = 256'hA59567F0600F79B4494445404A50B5504A69669664504A50B55B049A90570777;
defparam dpb_inst_4.INIT_RAM_0C = 256'h76615FBF69F7AF69F979A7797775A04B50B5504B6966966A504B50B550BA4B97;
defparam dpb_inst_4.INIT_RAM_0D = 256'hA04C50C5504C7477B77A504C50C550C64CB75AB5B66BF0600F0767A770777607;
defparam dpb_inst_4.INIT_RAM_0E = 256'h1111111F00F79F74F7876A8688665166780795073509595034579349977B7775;
defparam dpb_inst_4.INIT_RAM_0F = 256'hBA50A0BA777076779774504A50AA049A95765577077767766157606551111111;
defparam dpb_inst_4.INIT_RAM_10 = 256'hB0B9A5795556776507767766160F060001111111111111105577077559555450;
defparam dpb_inst_4.INIT_RAM_11 = 256'h076779774504A50AA049A97770767797775A04A50B04A77707677977A50BA50B;
defparam dpb_inst_4.INIT_RAM_12 = 256'h9BB5C55B5B66AF0600F446554565AA077760776615F0600F44540BA50A0BA777;
defparam dpb_inst_4.INIT_RAM_13 = 256'h7049504559095B505549B454B55B555590D5C0D550DC7477B77950BC50D550D6;
defparam dpb_inst_4.INIT_RAM_14 = 256'h006665550666060605555056556505F5BF74F5A7554745967774776878751778;
defparam dpb_inst_4.INIT_RAM_15 = 256'h000000000000000000000000000000000000000020F05025F55020F00F00025F;

DPB dpb_inst_5 (
    .DOA({dpb_inst_5_douta_w[11:0],douta[23:20]}),
    .DOB({dpb_inst_5_doutb_w[11:0],doutb[23:20]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[23:20]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[23:20]})
);

defparam dpb_inst_5.READ_MODE0 = 1'b1;
defparam dpb_inst_5.READ_MODE1 = 1'b1;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 4;
defparam dpb_inst_5.BIT_WIDTH_1 = 4;
defparam dpb_inst_5.BLK_SEL_0 = 3'b000;
defparam dpb_inst_5.BLK_SEL_1 = 3'b000;
defparam dpb_inst_5.RESET_MODE = "SYNC";
defparam dpb_inst_5.INIT_RAM_00 = 256'hC00048C0091DC0029100FD000140E20A0008C00FCCF1CE48F180000A08101D00;
defparam dpb_inst_5.INIT_RAM_01 = 256'hEDFF0E10000000010008C010F80809100000DE80C01E6080FAFFCFF0E10F140F;
defparam dpb_inst_5.INIT_RAM_02 = 256'h200E1E100042EBF20C048C048C048C048C02FEDC10FEDCBA9765105E1000C92F;
defparam dpb_inst_5.INIT_RAM_03 = 256'h8F518FA0C0D82983584185D8698F0986098589844983298210654329101D915F;
defparam dpb_inst_5.INIT_RAM_04 = 256'h10AF00E821E0FFCD0800F4EDCBA016C0C840C84000003290B100048C048C9411;
defparam dpb_inst_5.INIT_RAM_05 = 256'hE1404E3404D4DF000058400080ED000EDFF0E00EF0E10EE0000C048D15F01039;
defparam dpb_inst_5.INIT_RAM_06 = 256'h000404CF2002EE4F93E3DD4E91D1F000000000006543290C100FD0400002E808;
defparam dpb_inst_5.INIT_RAM_07 = 256'h00008000000040000000654329109D002905980000C48C048D4090009C050014;
defparam dpb_inst_5.INIT_RAM_08 = 256'hF010C020D020A000B001159291099006F000048C048C90050005C0100D8000C0;
defparam dpb_inst_5.INIT_RAM_09 = 256'h1000D0000D0000E8EFEFE0E0DE310E000C40000098764329815098810850F010;
defparam dpb_inst_5.INIT_RAM_0A = 256'hE310E0009ED3E10D800080048C04C048C50F3797A0001000D0009008F38D8A00;
defparam dpb_inst_5.INIT_RAM_0B = 256'hFE0FEF90D80D70F3696A000D00090005007F37D7A00D00090000900001CE0E0D;
defparam dpb_inst_5.INIT_RAM_0C = 256'h10F0D1E53ED3E53E1570F37F7A00050001000D005F35D5A0050001000D0E000B;
defparam dpb_inst_5.INIT_RAM_0D = 256'h040000000C002F72E2A0040000000C06000B6F0FD6FF90F8050DB1C6E00A4E03;
defparam dpb_inst_5.INIT_RAM_0E = 256'h4321980D00D7E57E9FCD06000CA0E06E604000400040000802080000F78F8A00;
defparam dpb_inst_5.INIT_RAM_0F = 256'h00080C006F3ED163F6A004000000800002B2F2EF0E0DE310E0C400000BA98765;
defparam dpb_inst_5.INIT_RAM_10 = 256'h0C0002B02EE2FEEC00DE310E000D0D8000C048C048C048C025A3FE153A5F000C;
defparam dpb_inst_5.INIT_RAM_11 = 256'hED163F6A008000400C00006F3ED163F6A0000000C00009E3FD193E9A00800040;
defparam dpb_inst_5.INIT_RAM_12 = 256'hF00504504D45490F8010099D0CBC5E0004E0310F0DD0D805A0000000C00006F3;
defparam dpb_inst_5.INIT_RAM_13 = 256'h600000000040000800000680F78B8A00040000000C008F78F8A0040000000C05;
defparam dpb_inst_5.INIT_RAM_14 = 256'h00011DCC0B11CB10F00000011C0100D7E57E95F549FAFD0733AFA0A0000D06D0;
defparam dpb_inst_5.INIT_RAM_15 = 256'h00000000000000000000000000000000000000000B1A0B0090000A10BDBBA005;

DPB dpb_inst_6 (
    .DOA({dpb_inst_6_douta_w[11:0],douta[27:24]}),
    .DOB({dpb_inst_6_doutb_w[11:0],doutb[27:24]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[27:24]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[27:24]})
);

defparam dpb_inst_6.READ_MODE0 = 1'b1;
defparam dpb_inst_6.READ_MODE1 = 1'b1;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 4;
defparam dpb_inst_6.BIT_WIDTH_1 = 4;
defparam dpb_inst_6.BLK_SEL_0 = 3'b000;
defparam dpb_inst_6.BLK_SEL_1 = 3'b000;
defparam dpb_inst_6.RESET_MODE = "SYNC";
defparam dpb_inst_6.INIT_RAM_00 = 256'h0001000E000A000100F00F00E00000000032200CDEE0EE6EE0E1E3EC322D0800;
defparam dpb_inst_6.INIT_RAM_01 = 256'h00FF0000C0C04C00F0100C10000C000F0C000000C00280C045000FF0000C0C0F;
defparam dpb_inst_6.INIT_RAM_02 = 256'h011222011000A0F05011112222333344444411111322222224444BBC00010030;
defparam dpb_inst_6.INIT_RAM_03 = 256'hE012E020203E14E15E16E16E17E028E119E10AE10BE10CE1001111100EEAEF70;
defparam dpb_inst_6.INIT_RAM_04 = 256'h000CC0000000006B3400222220011012111100000000332602C020001111C001;
defparam dpb_inst_6.INIT_RAM_05 = 256'h8088800000000F0000020000000000000FF00F00000000F00043333D06F3D030;
defparam dpb_inst_6.INIT_RAM_06 = 256'h000F064000001010000010100000100B00000000111110000E00000000008888;
defparam dpb_inst_6.INIT_RAM_07 = 256'h1000F0004000600040001111100E9240B00E42000210001117400004930200B3;
defparam dpb_inst_6.INIT_RAM_08 = 256'h800AA08AA00AA08AA0071F9100FA240B900020001111650F0048301009400020;
defparam dpb_inst_6.INIT_RAM_09 = 256'h000090001D01010100000200000002000650008011111132221D8EE799288088;
defparam dpb_inst_6.INIT_RAM_0A = 256'h0000E0009F41FD1C1103100000111222211F71010111B00040008000FB000011;
defparam dpb_inst_6.INIT_RAM_0B = 256'h00100011211A11F310101115000F0003001F7101011A000400018010100C2000;
defparam dpb_inst_6.INIT_RAM_0C = 256'h0040EEF91FD1F91F6111F31010111700010004001F7101011C00060009100010;
defparam dpb_inst_6.INIT_RAM_0D = 256'h10000A000D001FF1010115000F000211001010100100B1C11400000302005000;
defparam dpb_inst_6.INIT_RAM_0E = 256'h333222C90041F01F7F88111112010000011110210031110401111111FB101011;
defparam dpb_inst_6.INIT_RAM_0F = 256'h00090C0010100011030115000F01201011010100200000004065002001111133;
defparam dpb_inst_6.INIT_RAM_10 = 256'h1B0101011001C0002000000A000B1C110401111222233330110100011030111F;
defparam dpb_inst_6.INIT_RAM_11 = 256'h00011030112000C01F0101101000110301119000206000010000102011E00080;
defparam dpb_inst_6.INIT_RAM_12 = 256'h0011011110111A1A1190000000005020150000040E51611D0111D00060A00101;
defparam dpb_inst_6.INIT_RAM_13 = 256'h09010A0101B1110C11111111FF1010111800020005001F3101011D0007000A11;
defparam dpb_inst_6.INIT_RAM_14 = 256'h00E000000E000002F00660E000000011FD1FD101100000011100010111100001;
defparam dpb_inst_6.INIT_RAM_15 = 256'h00000000000000000000000000000000000000000060E000700000900900000B;

DPB dpb_inst_7 (
    .DOA({dpb_inst_7_douta_w[11:0],douta[31:28]}),
    .DOB({dpb_inst_7_doutb_w[11:0],doutb[31:28]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[31:28]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[31:28]})
);

defparam dpb_inst_7.READ_MODE0 = 1'b1;
defparam dpb_inst_7.READ_MODE1 = 1'b1;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 4;
defparam dpb_inst_7.BIT_WIDTH_1 = 4;
defparam dpb_inst_7.BLK_SEL_0 = 3'b000;
defparam dpb_inst_7.BLK_SEL_1 = 3'b000;
defparam dpb_inst_7.RESET_MODE = "SYNC";
defparam dpb_inst_7.INIT_RAM_00 = 256'h0600000F000F000000F00F06F00600006000000FFFF0FF4FF0F0F0FF000F0002;
defparam dpb_inst_7.INIT_RAM_01 = 256'h00FF000452520520F00005F00225200F052000225200305200000FF000450520;
defparam dpb_inst_7.INIT_RAM_02 = 256'h300000000003F0030000000000000000000300000000000000000FF502000E00;
defparam dpb_inst_7.INIT_RAM_03 = 256'h300C300400C30C30C30C30C30C300C300C300C300C300C30040000000FFEFDF0;
defparam dpb_inst_7.INIT_RAM_04 = 256'h000FF0000040040B0000000000000000000000000200000000F000000000F00C;
defparam dpb_inst_7.INIT_RAM_05 = 256'h0000000000000F03303238030000B00000F00000F00000F06000000F0B00F000;
defparam dpb_inst_7.INIT_RAM_06 = 256'h2007002000000000000000000000000200000000000000100F00000400030000;
defparam dpb_inst_7.INIT_RAM_07 = 256'h700060002000100020000000000FF902F00F9002000000000902D000902D0090;
defparam dpb_inst_7.INIT_RAM_08 = 256'h52C552C552C552C552CDDCC000FF802F600000000000802B000802C008020010;
defparam dpb_inst_7.INIT_RAM_09 = 256'h300020000200000000040000000011000100023000000000000FFE3E55D552C5;
defparam dpb_inst_7.INIT_RAM_0A = 256'h00010000FFF0FE0E0000000000000000000F00000000200020002004F0000000;
defparam dpb_inst_7.INIT_RAM_0B = 256'h000004F0F00E00F10000000100000001004F1000000100010000100000400000;
defparam dpb_inst_7.INIT_RAM_0C = 256'h01001EFE0FF0FF0FE040F00000000000000000004F0000000000000000000000;
defparam dpb_inst_7.INIT_RAM_0D = 256'h0700060006004F000000070006000700000000000004F0F00D00000000000020;
defparam dpb_inst_7.INIT_RAM_0E = 256'h000000FB00F0FF0FEFEE000000000000006000600060000600040000F0000000;
defparam dpb_inst_7.INIT_RAM_0F = 256'h0004040040040000000005000400500000000004000000011010023000000000;
defparam dpb_inst_7.INIT_RAM_10 = 256'h030000000000040400000011000E0E0000000000000000000400400000000004;
defparam dpb_inst_7.INIT_RAM_11 = 256'h4000000000300020020000400400000000003000303004004000000000300030;
defparam dpb_inst_7.INIT_RAM_12 = 256'h0000000000004F0F00D0040404000000000200100DE0E00D0000200020200400;
defparam dpb_inst_7.INIT_RAM_13 = 256'h000000000000000000000040F00000000100010001004F100000010001000100;
defparam dpb_inst_7.INIT_RAM_14 = 256'h00F000400F000000F00000F0000000F0FE0FB000040444000400000000000000;
defparam dpb_inst_7.INIT_RAM_15 = 256'h000000000000000000000000000000000000000004F4F400F00004F04F40400F;

endmodule //Gowin_DPB
