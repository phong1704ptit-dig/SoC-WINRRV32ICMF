// Created with Corsair v1.0.4

`ifndef __REGS_PWM_VH
`define __REGS_PWM_VH

`define PCSR_BASE_ADDR 0
`define PCSR_DATA_WIDTH 32
`define PCSR_ADDR_WIDTH 32

// TPWM_config - PWM configuration register
`define PCSR_TPWM_CONFIG_ADDR 32'h0
`define PCSR_TPWM_CONFIG_RESET 32'h0

// TPWM_config.EN - Enable PWM operation
`define PCSR_TPWM_CONFIG_EN_WIDTH 1
`define PCSR_TPWM_CONFIG_EN_LSB 0
`define PCSR_TPWM_CONFIG_EN_MASK 32'h0
`define PCSR_TPWM_CONFIG_EN_RESET 1'h0

// TPWM_config.SEL1 - Output selection for PWM1
`define PCSR_TPWM_CONFIG_SEL1_WIDTH 2
`define PCSR_TPWM_CONFIG_SEL1_LSB 1
`define PCSR_TPWM_CONFIG_SEL1_MASK 32'h0
`define PCSR_TPWM_CONFIG_SEL1_RESET 2'h0

// TPWM_config.SEL2 - Output selection for PWM2
`define PCSR_TPWM_CONFIG_SEL2_WIDTH 2
`define PCSR_TPWM_CONFIG_SEL2_LSB 3
`define PCSR_TPWM_CONFIG_SEL2_MASK 32'h0
`define PCSR_TPWM_CONFIG_SEL2_RESET 2'h0

// TPWM_config.RESERVED1 - Reserved for future use
`define PCSR_TPWM_CONFIG_RESERVED1_WIDTH 2
`define PCSR_TPWM_CONFIG_RESERVED1_LSB 5
`define PCSR_TPWM_CONFIG_RESERVED1_MASK 32'h0
`define PCSR_TPWM_CONFIG_RESERVED1_RESET 2'h0

// TPWM_config.SEL3 - Output selection for PWM3
`define PCSR_TPWM_CONFIG_SEL3_WIDTH 2
`define PCSR_TPWM_CONFIG_SEL3_LSB 7
`define PCSR_TPWM_CONFIG_SEL3_MASK 32'h0
`define PCSR_TPWM_CONFIG_SEL3_RESET 2'h0

// TPWM_config.SEL4 - Output selection for PWM4
`define PCSR_TPWM_CONFIG_SEL4_WIDTH 2
`define PCSR_TPWM_CONFIG_SEL4_LSB 9
`define PCSR_TPWM_CONFIG_SEL4_MASK 32'h0
`define PCSR_TPWM_CONFIG_SEL4_RESET 2'h0

// TPWM_config.NUM - Number of PWM signals selected
`define PCSR_TPWM_CONFIG_NUM_WIDTH 3
`define PCSR_TPWM_CONFIG_NUM_LSB 11
`define PCSR_TPWM_CONFIG_NUM_MASK 32'h0
`define PCSR_TPWM_CONFIG_NUM_RESET 3'h0

// TPWM_config.POL - Polarity of the PWM signal
`define PCSR_TPWM_CONFIG_POL_WIDTH 1
`define PCSR_TPWM_CONFIG_POL_LSB 14
`define PCSR_TPWM_CONFIG_POL_MASK 32'h0
`define PCSR_TPWM_CONFIG_POL_RESET 1'h0


// TPWM_prescaler - PWM clock divider
`define PCSR_TPWM_PRESCALER_ADDR 32'h4
`define PCSR_TPWM_PRESCALER_RESET 32'h1b

// TPWM_prescaler.DIV - Clock divider value for PWM
`define PCSR_TPWM_PRESCALER_DIV_WIDTH 32
`define PCSR_TPWM_PRESCALER_DIV_LSB 0
`define PCSR_TPWM_PRESCALER_DIV_MASK 32'h4
`define PCSR_TPWM_PRESCALER_DIV_RESET 32'h1b


// TPWM_period1 - PWM1 and PWM2 period register
`define PCSR_TPWM_PERIOD1_ADDR 32'h8
`define PCSR_TPWM_PERIOD1_RESET 32'hffffffff

// TPWM_period1.PER1 - Period value for PWM1
`define PCSR_TPWM_PERIOD1_PER1_WIDTH 16
`define PCSR_TPWM_PERIOD1_PER1_LSB 0
`define PCSR_TPWM_PERIOD1_PER1_MASK 32'h8
`define PCSR_TPWM_PERIOD1_PER1_RESET 16'hffff

// TPWM_period1.PER2 - Period value for PWM2
`define PCSR_TPWM_PERIOD1_PER2_WIDTH 16
`define PCSR_TPWM_PERIOD1_PER2_LSB 16
`define PCSR_TPWM_PERIOD1_PER2_MASK 32'h8
`define PCSR_TPWM_PERIOD1_PER2_RESET 16'hffff


// TPWM_period2 - PWM3 and PWM4 period register
`define PCSR_TPWM_PERIOD2_ADDR 32'hc
`define PCSR_TPWM_PERIOD2_RESET 32'hffffffff

// TPWM_period2.PER3 - Period value for PWM3
`define PCSR_TPWM_PERIOD2_PER3_WIDTH 16
`define PCSR_TPWM_PERIOD2_PER3_LSB 0
`define PCSR_TPWM_PERIOD2_PER3_MASK 32'hc
`define PCSR_TPWM_PERIOD2_PER3_RESET 16'hffff

// TPWM_period2.PER4 - Period value for PWM4
`define PCSR_TPWM_PERIOD2_PER4_WIDTH 16
`define PCSR_TPWM_PERIOD2_PER4_LSB 16
`define PCSR_TPWM_PERIOD2_PER4_MASK 32'hc
`define PCSR_TPWM_PERIOD2_PER4_RESET 16'hffff


// TPWM_compare1 - Compare values for PWM1 and PWM2
`define PCSR_TPWM_COMPARE1_ADDR 32'h10
`define PCSR_TPWM_COMPARE1_RESET 32'hffffffff

// TPWM_compare1.CP1 - Compare value for PWM1
`define PCSR_TPWM_COMPARE1_CP1_WIDTH 16
`define PCSR_TPWM_COMPARE1_CP1_LSB 0
`define PCSR_TPWM_COMPARE1_CP1_MASK 32'h10
`define PCSR_TPWM_COMPARE1_CP1_RESET 16'hffff

// TPWM_compare1.CP2 - Compare value for PWM2
`define PCSR_TPWM_COMPARE1_CP2_WIDTH 16
`define PCSR_TPWM_COMPARE1_CP2_LSB 16
`define PCSR_TPWM_COMPARE1_CP2_MASK 32'h10
`define PCSR_TPWM_COMPARE1_CP2_RESET 16'hffff


// TPWM_compare2 - Compare values for PWM3 and PWM4
`define PCSR_TPWM_COMPARE2_ADDR 32'h14
`define PCSR_TPWM_COMPARE2_RESET 32'hffffffff

// TPWM_compare2.CP3 - Compare value for PWM3
`define PCSR_TPWM_COMPARE2_CP3_WIDTH 16
`define PCSR_TPWM_COMPARE2_CP3_LSB 0
`define PCSR_TPWM_COMPARE2_CP3_MASK 32'h14
`define PCSR_TPWM_COMPARE2_CP3_RESET 16'hffff

// TPWM_compare2.CP4 - Compare value for PWM4
`define PCSR_TPWM_COMPARE2_CP4_WIDTH 16
`define PCSR_TPWM_COMPARE2_CP4_LSB 16
`define PCSR_TPWM_COMPARE2_CP4_MASK 32'h14
`define PCSR_TPWM_COMPARE2_CP4_RESET 16'hffff


// TPWM_counter1 - PWM counters for PWM1 and PWM2
`define PCSR_TPWM_COUNTER1_ADDR 32'h18
`define PCSR_TPWM_COUNTER1_RESET 32'h0

// TPWM_counter1.CNT1 - Current counter value for PWM1
`define PCSR_TPWM_COUNTER1_CNT1_WIDTH 16
`define PCSR_TPWM_COUNTER1_CNT1_LSB 0
`define PCSR_TPWM_COUNTER1_CNT1_MASK 32'h18
`define PCSR_TPWM_COUNTER1_CNT1_RESET 16'h0

// TPWM_counter1.CNT2 - Current counter value for PWM2
`define PCSR_TPWM_COUNTER1_CNT2_WIDTH 16
`define PCSR_TPWM_COUNTER1_CNT2_LSB 16
`define PCSR_TPWM_COUNTER1_CNT2_MASK 32'h18
`define PCSR_TPWM_COUNTER1_CNT2_RESET 16'h0


// TPWM_counter2 - PWM counters for PWM3 and PWM4
`define PCSR_TPWM_COUNTER2_ADDR 32'h1c
`define PCSR_TPWM_COUNTER2_RESET 32'h0

// TPWM_counter2.CNT3 - Current counter value for PWM3
`define PCSR_TPWM_COUNTER2_CNT3_WIDTH 16
`define PCSR_TPWM_COUNTER2_CNT3_LSB 0
`define PCSR_TPWM_COUNTER2_CNT3_MASK 32'h1c
`define PCSR_TPWM_COUNTER2_CNT3_RESET 16'h0

// TPWM_counter2.CNT4 - Current counter value for PWM4
`define PCSR_TPWM_COUNTER2_CNT4_WIDTH 16
`define PCSR_TPWM_COUNTER2_CNT4_LSB 16
`define PCSR_TPWM_COUNTER2_CNT4_MASK 32'h1c
`define PCSR_TPWM_COUNTER2_CNT4_RESET 16'h0


`endif // __REGS_PWM_VH